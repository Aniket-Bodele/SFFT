`timescale 1ns/1ps
`include"sfft.v"
module sfft_test ;
reg [11:0] in0_r,in0_i,in1_r,in1_i,in2_r,in2_i,in3_r,in3_i,in4_r,in4_i,in5_r,in5_i,in6_r,in6_i,
            in7_r,in7_i,in8_r,in8_i,in9_r,in9_i,in10_r,in10_i,in11_r,in11_i,in12_r,in12_i,in13_r,in13_i,
            in14_r,in14_i,in15_r,in15_i,in16_r,in16_i,in17_r,in17_i,in18_r,in18_i,in19_r,in19_i,in20_r,in20_i,
            in21_r,in21_i,in22_r,in22_i,in23_r,in23_i,in24_r,in24_i,in25_r,in25_i,in26_r,in26_i,in27_r,in27_i,
            in28_r,in28_i,in29_r,in29_i,in30_r,in30_i,in31_r,in31_i,in32_r,in32_i,in33_r,in33_i,in34_r,in34_i,
            in35_r,in35_i,in36_r,in36_i,in37_r,in37_i,in38_r,in38_i,in39_r,in39_i,in40_r,in40_i,in41_r,in41_i,
            in42_r,in42_i,in43_r,in43_i,in44_r,in44_i,in45_r,in45_i,in46_r,in46_i,in47_r,in47_i,in48_r,in48_i,
            in49_r,in49_i,in50_r,in50_i,in51_r,in51_i,in52_r,in52_i,in53_r,in53_i,in54_r,in54_i,in55_r,in55_i,
            in56_r,in56_i,in57_r,in57_i,in58_r,in58_i,in59_r,in59_i,in60_r,in60_i,in61_r,in61_i,
            in62_r,in62_i,in63_r,in63_i; 
reg clk;
wire [11:0] y0_r,y0_i,y1_r,y1_i,y2_r,y2_i,y3_r,y3_i,y4_r,y4_i,y5_r,y5_i,y6_r,y6_i,y7_r,y7_i,y8_r,y8_i,y9_r,y9_i,
y10_r,y10_i,y11_r,y11_i,y12_r,y12_i,y13_r,y13_i,y14_r,y14_i,y15_r,y15_i,y16_r,y16_i,y17_r,y17_i,y18_r,y18_i,y19_r,y19_i,y20_r,y20_i,y21_r,y21_i,
y22_r,y22_i,y23_r,y23_i,y24_r,y24_i,y25_r,y25_i,y26_r,y26_i,y27_r,y27_i,y28_r,y28_i,y29_r,y29_i,y30_r,y30_i,y31_r,y31_i,y32_r,y32_i,y33_r,y33_i,y34_r,y34_i,y35_r,y35_i,y36_r,y36_i,y37_r,y37_i,y38_r,y38_i,y39_r,y39_i,
y40_r,y40_i,y41_r,y41_i,y42_r,y42_i,y43_r,y43_i,y44_r,y44_i,y45_r,y45_i,y46_r,y46_i,y47_r,y47_i,y48_r,y48_i,y49_r,y49_i,y50_r,y50_i,y51_r,y51_i,
y52_r,y52_i,y53_r,y53_i,y54_r,y54_i,y55_r,y55_i,y56_r,y56_i,y57_r,y57_i,y58_r,y58_i,y59_r,y59_i,y60_r,y60_i,y61_r,y61_i,y62_r,y62_i,y63_r,y63_i;


SFFT SFFT (in0_r,in0_i,y0_r,y0_i,
in1_r,in1_i,y1_r,y1_i,
in2_r,in2_i,y2_r,y2_i,
in3_r,in3_i,y3_r,y3_i,
in4_r,in4_i,y4_r,y4_i,
in5_r,in5_i,y5_r,y5_i,
in6_r,in6_i,y6_r,y6_i,
in7_r,in7_i,y7_r,y7_i,
in8_r,in8_i,y8_r,y8_i,
in9_r,in9_i,y9_r,y9_i,
in10_r,in10_i,y10_r,y10_i,
in11_r,in11_i,y11_r,y11_i,
in12_r,in12_i,y12_r,y12_i,
in13_r,in13_i,y13_r,y13_i,
in14_r,in14_i,y14_r,y14_i,
in15_r,in15_i,y15_r,y15_i,
in16_r,in16_i,y16_r,y16_i,
in17_r,in17_i,y17_r,y17_i,
in18_r,in18_i,y18_r,y18_i,
in19_r,in19_i,y19_r,y19_i,
in20_r,in20_i,y20_r,y20_i,
in21_r,in21_i,y21_r,y21_i,
in22_r,in22_i,y22_r,y22_i,
in23_r,in23_i,y23_r,y23_i,
in24_r,in24_i,y24_r,y24_i,
in25_r,in25_i,y25_r,y25_i,
in26_r,in26_i,y26_r,y26_i,
in27_r,in27_i,y27_r,y27_i,
in28_r,in28_i,y28_r,y28_i,
in29_r,in29_i,y29_r,y29_i,
in30_r,in30_i,y30_r,y30_i,
in31_r,in31_i,y31_r,y31_i,
in32_r,in32_i,y32_r,y32_i,
in33_r,in33_i,y33_r,y33_i,
in34_r,in34_i,y34_r,y34_i,
in35_r,in35_i,y35_r,y35_i,
in36_r,in36_i,y36_r,y36_i,
in37_r,in37_i,y37_r,y37_i,
in38_r,in38_i,y38_r,y38_i,
in39_r,in39_i,y39_r,y39_i,
in40_r,in40_i,y40_r,y40_i,
in41_r,in41_i,y41_r,y41_i,
in42_r,in42_i,y42_r,y42_i,
in43_r,in43_i,y43_r,y43_i,
in44_r,in44_i,y44_r,y44_i,
in45_r,in45_i,y45_r,y45_i,
in46_r,in46_i,y46_r,y46_i,
in47_r,in47_i,y47_r,y47_i,
in48_r,in48_i,y48_r,y48_i,
in49_r,in49_i,y49_r,y49_i,
in50_r,in50_i,y50_r,y50_i,
in51_r,in51_i,y51_r,y51_i,
in52_r,in52_i,y52_r,y52_i,
in53_r,in53_i,y53_r,y53_i,
in54_r,in54_i,y54_r,y54_i,
in55_r,in55_i,y55_r,y55_i,
in56_r,in56_i,y56_r,y56_i,
in57_r,in57_i,y57_r,y57_i,
in58_r,in58_i,y58_r,y58_i,
in59_r,in59_i,y59_r,y59_i,
in60_r,in60_i,y60_r,y60_i,
in61_r,in61_i,y61_r,y61_i,
in62_r,in62_i,y62_r,y62_i,
in63_r,in63_i,y63_r,y63_i,clk);



initial
begin
    clk=1'b0;
    #1000 $finish;
end
always #5 clk=~clk;  
initial
begin
    in0_r=12'b000000000000; 
    in1_r=12'b000000100000;
    in2_r=12'b000010000000;
    in3_r=12'b000001000000;
    in4_r=12'b000000010000;
    in5_r=12'b000001100000;
    in6_r=12'b000000110000;
    in7_r=12'b000001010000;
    in8_r=12'b000001010000;
    in9_r=12'b000001000000;
   in10_r=12'b000000110000;
   in11_r=12'b000000010000;
   in12_r=12'b000000100000;
   in13_r=12'b000010000000;
   in14_r=12'b000001110000;
   in15_r=12'b000010010000;
   in16_r=12'b000000010000;
   in17_r=12'b000001110000;
   in18_r=12'b000001010000;
   in19_r=12'b000001000000;
   in20_r=12'b000000110000;
   in21_r=12'b000000100000;
   in22_r=12'b000010000000;
   in23_r=12'b000001100000;
   in24_r=12'b000000000000;
   in25_r=12'b000010010000;
   in26_r=12'b000000010000;
   in27_r=12'b000000010000;
   in28_r=12'b000001010000;
   in29_r=12'b000001110000;
   in30_r=12'b000010000000;
   in31_r=12'b000001000000;
   in32_r=12'b000001000000;
   in33_r=12'b000000000000;
   in34_r=12'b000000000000;
   in35_r=12'b000000000000;
   in36_r=12'b000010010000;
   in37_r=12'b000000010000;
   in38_r=12'b000000100000;
   in39_r=12'b000000110000;
   in40_r=12'b000000110000;
   in41_r=12'b000000100000;
   in42_r=12'b000000010000;
   in43_r=12'b000010010000;
   in44_r=12'b000000000000;
   in45_r=12'b000000000000;
   in46_r=12'b000000000000;
   in47_r=12'b000000000000;
   in48_r=12'b000000100000;
   in49_r=12'b000000010000;
   in50_r=12'b000001000000;
   in51_r=12'b000001000000;
   in52_r=12'b000000110000;
   in53_r=12'b000010010000;
   in54_r=12'b000000000000;
   in55_r=12'b000000010000;
   in56_r=12'b000000010000;
   in57_r=12'b000000010000;
   in58_r=12'b000000010000;
   in59_r=12'b000000100000;
   in60_r=12'b000000100000;
   in61_r=12'b000000010000;
   in62_r=12'b000000010000;
   in63_r=12'b000000010000;

 in0_i=12'b000000000000;
 in1_i=12'b000000000000;
 in2_i=12'b000000000000;
 in3_i=12'b000000000000;
 in4_i=12'b000000000000;
 in5_i=12'b000000000000;
 in6_i=12'b000000000000;
 in7_i=12'b000000000000;
 in8_i=12'b000000000000;
 in9_i=12'b000000000000;
in10_i=12'b000000000000;
in11_i=12'b000000000000;
in12_i=12'b000000000000;
in13_i=12'b000000000000;
in14_i=12'b000000000000;
in15_i=12'b000000000000;
in16_i=12'b000000000000;
in17_i=12'b000000000000;
in18_i=12'b000000000000;
in19_i=12'b000000000000;
in20_i=12'b000000000000;
in21_i=12'b000000000000;
in22_i=12'b000000000000;
in23_i=12'b000000000000;
in24_i=12'b000000000000;
in25_i=12'b000000000000;
in26_i=12'b000000000000;
in27_i=12'b000000000000;
in28_i=12'b000000000000;
in29_i=12'b000000000000;
in30_i=12'b000000000000;
in31_i=12'b000000000000;
in32_i=12'b000000000000;
in33_i=12'b000000000000;
in34_i=12'b000000000000;
in35_i=12'b000000000000;
in36_i=12'b000000000000;
in37_i=12'b000000000000;
in38_i=12'b000000000000;
in39_i=12'b000000000000;
in40_i=12'b000000000000;
in41_i=12'b000000000000;
in42_i=12'b000000000000;
in43_i=12'b000000000000;
in44_i=12'b000000000000;
in45_i=12'b000000000000;
in46_i=12'b000000000000;
in47_i=12'b000000000000;
in48_i=12'b000000000000;
in49_i=12'b000000000000;
in50_i=12'b000000000000;
in51_i=12'b000000000000;
in52_i=12'b000000000000;
in53_i=12'b000000000000;
in54_i=12'b000000000000;
in55_i=12'b000000000000;
in56_i=12'b000000000000;
in57_i=12'b000000000000;
in58_i=12'b000000000000;
in59_i=12'b000000000000;
in60_i=12'b000000000000;
in61_i=12'b000000000000;
in62_i=12'b000000000000;
in63_i=12'b000000000000;
end
initial
begin
    
    $dumpfile("sfft.vcd");$dumpvars(0,sfft_test);
end
    
endmodule